library verilog;
use verilog.vl_types.all;
entity alu_control is
    port(
        opcode          : in     vl_logic_vector(6 downto 0);
        funct3          : in     vl_logic_vector(2 downto 0);
        funct7          : in     vl_logic_vector(6 downto 0);
        alu_ctrl        : out    vl_logic_vector(3 downto 0)
    );
end alu_control;
